module decoder
{
    iRst,
    imData,
    imData_Ready,
    oCode,
    oCode_Ready

};


// ==== I/O, Reg, Wire Declaration ======================================
input       [7:0]               imData;
input                           imData_Ready;



output      [7:0]               oCode;
output                          oCode_Ready;
                

// ==== Structural Design ==============================




endmodule